
module tan_lut (
    input [6-1:0] num,
    output reg [25-1:0] atan
);

wire signed [25-1:0] atan_table [0:22];

assign atan_table[0] = 25'b0011001001000011111101101;
assign atan_table[1] = 25'b0001110110101100011001110;
assign atan_table[2] = 25'b0000111110101101101110101;
assign atan_table[3] = 25'b0000011111110101011011101;
assign atan_table[4] = 25'b0000001111111110101010110;
assign atan_table[5] = 25'b0000000111111111110101010;
assign atan_table[6] = 25'b0000000011111111111110101;
assign atan_table[7] = 25'b0000000001111111111111110;
assign atan_table[8] = 25'b0000000000111111111111111;
assign atan_table[9] = 25'b0000000000011111111111111;
assign atan_table[10] = 25'b0000000000001111111111111;
assign atan_table[11] = 25'b0000000000000111111111111;
assign atan_table[12] = 25'b0000000000000011111111111;
assign atan_table[13] = 25'b0000000000000001111111111;
assign atan_table[14] = 25'b0000000000000000111111111;
assign atan_table[15] = 25'b0000000000000000011111111;
assign atan_table[16] = 25'b0000000000000000001111111;
assign atan_table[17] = 25'b0000000000000000000111111;
assign atan_table[18] = 25'b0000000000000000000011111;
assign atan_table[19] = 25'b0000000000000000000001111;
assign atan_table[20] = 25'b0000000000000000000000111;
assign atan_table[21] = 25'b0000000000000000000000011;
assign atan_table[22] = 25'b0000000000000000000000001;

always @(*) begin
    atan = atan_table[num];
end

endmodule